// arbiter.vh

`define IDLE 2'b00
`define GNT2 2'b01
`define GNT1 2'b10
`define GNT0 2'b11